--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   16:11:50 07/26/2022
-- Design Name:   
-- Module Name:   C:/Users/Hilary Calva Camacho/Desktop/PROYECTOS VHDL/GeneracionComponentes/TB_ProyectoContador.vhd
-- Project Name:  GeneracionComponentes
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: ProyectoContador
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
ENTITY TB_ProyectoContador IS
END TB_ProyectoContador;
 
ARCHITECTURE behavior OF TB_ProyectoContador IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT ProyectoContador
    PORT(
         clk : IN  std_logic;
         rst : IN  std_logic;
         display : OUT  std_logic_vector(6 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal clk : std_logic := '0';
   signal rst : std_logic := '0';

 	--Outputs
   signal display : std_logic_vector(6 downto 0);

   -- Clock period definitions
   constant clk_period : time := 10 ns;
 
BEGIN


 
	-- Instantiate the Unit Under Test (UUT)
   uut: ProyectoContador PORT MAP (
          clk => clk,
          rst => rst,
          display => display
        );

   -- Clock process definitions
   clk_process :process
   begin
		clk <= '0';
		wait for clk_period/2;
		clk <= '1';
		wait for clk_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		

      wait for clk_period*10;
		rst <= '0';
		wait for clk_period*10;
		rst <= '1';

      -- insert stimulus here 

      wait;
   end process;

END;
